module top_module ( input a, input b, output out );
    mod_a M(a,b,out);
endmodule
